package apb_pkg;
	
    `include "sequence_item.sv"
	`include "sequence.sv"
	`include "apb_sequencer.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "agent.sv"
	`include "predictor.sv"
	`include "scoreboard.sv"
	`include "environment.sv"
	//`include "write_test.sv"
//	`include "apb_read_test.sv"
//	`include "apb_random_write_read.sv"
//	`include "apb_pslverr_check.sv"
	`include "test.sv"
	event e1;
endpackage : apb_pkg
